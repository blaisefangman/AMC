magic
tech scmos
timestamp 1614220983
<< nwell >>
rect -4 210 36 248
rect -4 114 36 187
rect -4 0 36 54
<< pwell >>
rect -4 187 36 210
rect -4 54 36 114
<< ntransistor >>
rect 7 195 9 199
rect 15 195 17 199
rect 23 195 25 199
rect 15 89 17 102
rect 23 89 25 102
rect 7 69 9 73
rect 15 60 17 73
rect 23 60 25 73
<< ptransistor >>
rect 14 224 16 231
rect 22 224 24 231
rect 7 174 9 181
rect 15 174 17 181
rect 23 174 25 181
rect 15 120 17 146
rect 23 120 25 146
rect 7 41 9 48
rect 15 22 17 48
rect 23 22 25 48
<< ndiffusion >>
rect 6 195 7 199
rect 9 195 15 199
rect 17 195 18 199
rect 22 195 23 199
rect 25 195 26 199
rect 14 89 15 102
rect 17 89 18 102
rect 22 89 23 102
rect 25 89 26 102
rect 6 69 7 73
rect 9 69 10 73
rect 14 60 15 73
rect 17 60 18 73
rect 22 60 23 73
rect 25 60 26 73
<< pdiffusion >>
rect 13 224 14 231
rect 16 224 17 231
rect 21 224 22 231
rect 24 224 25 231
rect 6 174 7 181
rect 9 174 10 181
rect 14 174 15 181
rect 17 174 18 181
rect 22 174 23 181
rect 25 174 26 181
rect 14 120 15 146
rect 17 120 18 146
rect 22 120 23 146
rect 25 120 26 146
rect 6 41 7 48
rect 9 41 10 48
rect 14 22 15 48
rect 17 22 18 48
rect 22 22 23 48
rect 25 22 26 48
<< ndcontact >>
rect 2 195 6 199
rect 18 195 22 199
rect 26 195 30 199
rect 10 89 14 102
rect 18 89 22 102
rect 26 89 30 102
rect 2 69 6 73
rect 10 60 14 73
rect 18 60 22 73
rect 26 60 30 73
<< pdcontact >>
rect 9 224 13 231
rect 17 224 21 231
rect 25 224 29 231
rect 2 174 6 181
rect 10 174 14 181
rect 18 174 22 181
rect 26 174 30 181
rect 10 120 14 146
rect 18 120 22 146
rect 26 120 30 146
rect 2 41 6 48
rect 10 22 14 48
rect 18 22 22 48
rect 26 22 30 48
<< psubstratepcontact >>
rect 22 203 26 207
rect 26 81 30 85
<< nsubstratencontact >>
rect 17 216 21 220
rect 2 146 6 150
rect 14 14 18 18
<< polysilicon >>
rect 14 233 24 235
rect 14 231 16 233
rect 22 231 24 233
rect 14 222 16 224
rect 22 222 24 224
rect 6 216 9 221
rect 7 199 9 216
rect 16 208 17 210
rect 15 199 17 208
rect 23 199 25 201
rect 7 181 9 195
rect 15 181 17 195
rect 23 192 25 195
rect 24 188 25 192
rect 23 181 25 188
rect 7 172 9 174
rect 15 172 17 174
rect 7 110 9 165
rect 15 146 17 148
rect 23 146 25 174
rect 15 102 17 120
rect 23 118 25 120
rect 23 116 33 118
rect 24 106 25 110
rect 23 102 25 106
rect 15 80 17 89
rect 7 78 17 80
rect 7 73 9 78
rect 15 73 17 75
rect 23 73 25 89
rect 7 48 9 69
rect 15 56 17 60
rect 23 58 25 60
rect 31 52 33 116
rect 15 48 17 52
rect 23 50 33 52
rect 23 48 25 50
rect 7 11 9 41
rect 15 20 17 22
rect 23 20 25 22
rect 7 9 11 11
<< polycontact >>
rect 17 235 21 239
rect 2 216 6 220
rect 12 208 16 212
rect 20 188 24 192
rect 9 161 13 165
rect 7 106 11 110
rect 20 106 24 110
rect 13 52 17 56
rect 11 7 15 11
<< metal1 >>
rect 0 239 34 241
rect 0 238 17 239
rect 21 238 34 239
rect 0 212 34 213
rect 0 210 12 212
rect 16 210 34 212
rect 0 202 2 205
rect 19 205 22 206
rect 6 202 22 205
rect 18 199 22 202
rect 2 191 6 195
rect 2 188 20 191
rect 10 181 14 188
rect 27 181 30 195
rect 2 171 6 174
rect 18 171 22 174
rect 2 168 22 171
rect 26 165 30 174
rect 13 161 30 165
rect 14 154 30 157
rect 6 146 10 150
rect 26 146 30 154
rect 11 106 20 110
rect 27 102 30 120
rect 10 85 14 89
rect 0 81 10 85
rect 14 81 26 85
rect 30 81 34 85
rect 2 56 6 69
rect 2 52 13 56
rect 2 48 6 52
rect 26 48 30 60
rect 10 18 14 22
rect 0 14 14 18
rect 22 14 34 18
<< m2contact >>
rect 9 231 13 235
rect 25 231 29 235
rect 2 220 6 224
rect 17 220 21 224
rect 2 202 6 206
rect 18 181 22 185
rect 10 154 14 158
rect 10 146 14 150
rect 10 81 14 85
rect 10 73 14 77
rect 26 73 30 77
rect 18 14 22 18
rect 15 7 19 11
rect 5 0 9 4
<< metal2 >>
rect 9 235 12 248
rect 10 211 13 231
rect 22 231 25 248
rect 22 227 30 231
rect 6 202 7 205
rect 4 85 7 202
rect 10 158 14 211
rect 18 185 21 220
rect 18 150 21 181
rect 14 146 21 150
rect 4 81 10 85
rect 10 77 14 81
rect 18 18 21 146
rect 26 77 30 227
rect 4 5 5 9
rect 9 5 10 9
rect 4 4 10 5
rect 4 0 5 4
rect 9 0 10 4
rect 15 0 18 7
<< m3contact >>
rect 3 224 7 228
rect 5 5 9 9
<< metal3 >>
rect 2 228 10 229
rect 2 224 3 228
rect 7 224 10 228
rect 2 223 10 224
rect 4 9 10 223
rect 4 5 5 9
rect 9 5 10 9
rect 4 0 10 5
<< m3p >>
rect 0 0 34 248
<< labels >>
rlabel metal1 34 14 34 14 7 vdd
rlabel metal1 34 81 34 81 7 gnd
rlabel metal1 34 210 34 210 1 en
rlabel metal1 34 238 34 238 7 pchg
rlabel metal2 28 170 28 170 1 en1
rlabel polycontact 24 189 24 189 1 en_bar
rlabel metal2 9 248 9 248 5 br
rlabel metal2 22 248 22 248 5 bl
rlabel metal2 15 0 15 0 1 din
rlabel metal3 4 0 4 0 1 bm
<< end >>
