magic
tech scmos
timestamp 1614052413
<< nwell >>
rect 0 0 25 51
<< pwell >>
rect 25 0 50 51
<< ntransistor >>
rect 31 20 39 22
rect 31 12 39 14
<< ptransistor >>
rect 11 36 19 38
rect 11 28 19 30
rect 11 20 19 22
rect 11 12 19 14
<< ndiffusion >>
rect 31 23 33 27
rect 37 23 39 27
rect 31 22 39 23
rect 31 19 39 20
rect 31 15 33 19
rect 37 15 39 19
rect 31 14 39 15
rect 31 11 39 12
rect 31 7 33 11
rect 37 7 39 11
<< pdiffusion >>
rect 11 39 13 43
rect 17 39 19 43
rect 11 38 19 39
rect 11 35 19 36
rect 11 31 13 35
rect 17 31 19 35
rect 11 30 19 31
rect 11 27 19 28
rect 11 23 13 27
rect 17 23 19 27
rect 11 22 19 23
rect 11 19 19 20
rect 11 15 13 19
rect 17 15 19 19
rect 11 14 19 15
rect 11 11 19 12
rect 11 7 13 11
rect 17 7 19 11
<< ndcontact >>
rect 33 23 37 27
rect 33 15 37 19
rect 33 7 37 11
<< pdcontact >>
rect 13 39 17 43
rect 13 31 17 35
rect 13 23 17 27
rect 13 15 17 19
rect 13 7 17 11
<< psubstratepcontact >>
rect 33 40 37 44
<< nsubstratencontact >>
rect 3 38 7 42
<< polysilicon >>
rect 9 36 11 38
rect 19 37 31 38
rect 19 36 42 37
rect 29 35 42 36
rect 9 28 11 30
rect 19 29 46 30
rect 19 28 42 29
rect 9 20 11 22
rect 19 20 24 22
rect 28 20 31 22
rect 39 20 41 22
rect 5 12 11 14
rect 19 12 31 14
rect 39 12 41 14
<< polycontact >>
rect 42 33 46 37
rect 42 25 46 29
rect 24 18 28 22
rect 5 8 9 12
<< metal1 >>
rect 0 50 50 51
rect 0 47 9 50
rect 3 42 6 47
rect 13 47 50 50
rect 0 32 13 35
rect 17 31 37 34
rect 46 34 50 37
rect 33 27 37 31
rect 46 25 50 28
rect 0 9 5 12
rect 24 11 27 18
rect 17 7 33 11
rect 0 0 40 4
rect 44 0 50 4
<< m2contact >>
rect 9 46 13 50
rect 17 39 21 43
rect 37 40 41 44
rect 17 23 21 27
rect 9 15 13 19
rect 37 15 41 19
rect 40 0 44 4
<< metal2 >>
rect 9 19 12 46
rect 21 23 24 43
rect 41 4 44 44
<< m3p >>
rect 0 0 50 51
<< labels >>
rlabel metal1 0 49 0 49 8 vdd
rlabel metal1 0 2 0 2 6 gnd
rlabel metal1 0 32 0 32 3 dr
rlabel metal1 0 9 0 9 3 sen
rlabel metal1 50 25 50 25 7 bl
rlabel metal1 50 34 50 34 7 br
<< end >>
