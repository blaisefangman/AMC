magic
tech scmos
timestamp 1615313102
<< nwell >>
rect -2 254 19 344
rect -2 92 17 254
rect -2 0 19 92
<< pwell >>
rect 19 254 36 344
rect 17 92 36 254
rect 19 0 36 92
<< ntransistor >>
rect 26 293 30 313
rect 26 283 30 287
rect 26 267 30 269
rect 23 228 30 230
rect 23 220 30 222
rect 23 211 30 213
rect 23 202 30 204
rect 23 151 30 153
rect 23 142 30 144
rect 23 133 30 135
rect 23 117 30 119
rect 26 79 30 81
rect 26 65 30 67
rect 26 47 30 51
rect 26 21 30 41
<< ptransistor >>
rect 5 293 13 313
rect 5 283 13 287
rect 5 267 13 269
rect 5 245 11 247
rect 5 220 11 222
rect 5 202 11 204
rect 5 151 11 153
rect 5 133 11 135
rect 5 100 11 102
rect 5 79 13 81
rect 5 65 13 67
rect 5 47 13 51
rect 5 21 13 41
<< ndiffusion >>
rect 26 313 30 314
rect 26 292 30 293
rect 29 288 30 292
rect 26 287 30 288
rect 26 282 30 283
rect 29 278 30 282
rect 29 270 30 274
rect 26 269 30 270
rect 26 266 30 267
rect 27 237 30 241
rect 23 230 30 237
rect 23 222 30 228
rect 23 213 30 220
rect 23 204 30 211
rect 23 201 30 202
rect 23 197 26 201
rect 23 154 26 158
rect 23 153 30 154
rect 23 144 30 151
rect 23 135 30 142
rect 23 119 30 133
rect 23 110 30 117
rect 27 106 30 110
rect 29 82 30 86
rect 26 81 30 82
rect 26 72 30 79
rect 26 67 30 68
rect 26 64 30 65
rect 29 60 30 64
rect 29 52 30 56
rect 26 51 30 52
rect 26 41 30 47
rect 26 20 30 21
<< pdiffusion >>
rect 9 314 13 318
rect 5 313 13 314
rect 5 292 13 293
rect 9 288 13 292
rect 5 287 13 288
rect 5 282 13 283
rect 9 278 13 282
rect 9 270 13 274
rect 5 269 13 270
rect 5 266 13 267
rect 9 262 13 266
rect 9 250 11 254
rect 5 247 11 250
rect 5 244 11 245
rect 9 240 11 244
rect 9 223 11 227
rect 5 222 11 223
rect 5 204 11 220
rect 5 201 11 202
rect 9 197 11 201
rect 9 154 11 158
rect 5 153 11 154
rect 5 135 11 151
rect 5 132 11 133
rect 9 128 11 132
rect 9 103 11 107
rect 5 102 11 103
rect 5 97 11 100
rect 9 93 11 97
rect 9 82 13 86
rect 5 81 13 82
rect 5 72 13 79
rect 9 68 13 72
rect 5 67 13 68
rect 5 64 13 65
rect 9 60 13 64
rect 9 52 13 56
rect 5 51 13 52
rect 5 41 13 47
rect 5 20 13 21
rect 9 16 13 20
<< ndcontact >>
rect 26 314 30 318
rect 25 288 29 292
rect 25 278 29 282
rect 25 270 29 274
rect 26 262 30 266
rect 23 237 27 241
rect 26 197 30 201
rect 26 154 30 158
rect 23 106 27 110
rect 25 82 29 86
rect 26 68 30 72
rect 25 60 29 64
rect 25 52 29 56
rect 26 16 30 20
<< pdcontact >>
rect 5 314 9 318
rect 5 288 9 292
rect 5 278 9 282
rect 5 270 9 274
rect 5 262 9 266
rect 5 250 9 254
rect 5 240 9 244
rect 5 223 9 227
rect 5 197 9 201
rect 5 154 9 158
rect 5 128 9 132
rect 5 103 9 107
rect 5 93 9 97
rect 5 82 9 86
rect 5 68 9 72
rect 5 60 9 64
rect 5 52 9 56
rect 5 16 9 20
<< psubstratepcontact >>
rect 26 323 30 327
rect 26 4 30 8
<< nsubstratencontact >>
rect 5 323 9 327
rect 5 4 9 8
<< polysilicon >>
rect 2 293 5 313
rect 13 312 16 313
rect 13 308 14 312
rect 13 293 16 308
rect 24 305 26 313
rect 25 301 26 305
rect 24 293 26 301
rect 30 293 32 313
rect 3 283 5 287
rect 13 284 16 287
rect 20 284 26 287
rect 13 283 26 284
rect 30 283 32 287
rect 3 267 5 269
rect 13 268 26 269
rect 13 267 16 268
rect 20 267 26 268
rect 30 267 32 269
rect 3 245 5 247
rect 11 245 13 247
rect 21 228 23 230
rect 30 228 32 230
rect 3 220 5 222
rect 11 220 23 222
rect 30 220 32 222
rect 15 209 16 213
rect 20 211 23 213
rect 30 211 32 213
rect 3 202 5 204
rect 11 202 23 204
rect 30 202 32 204
rect 3 151 5 153
rect 11 151 23 153
rect 30 151 32 153
rect 21 142 23 144
rect 30 142 32 144
rect 3 133 5 135
rect 11 133 23 135
rect 30 133 32 135
rect 17 117 23 119
rect 30 117 32 119
rect 3 100 5 102
rect 11 100 13 102
rect 3 79 5 81
rect 13 79 18 81
rect 22 79 26 81
rect 30 79 32 81
rect 3 65 5 67
rect 13 66 16 67
rect 20 66 26 67
rect 13 65 26 66
rect 30 65 32 67
rect 3 47 5 51
rect 13 50 26 51
rect 13 47 16 50
rect 20 47 26 50
rect 30 47 32 51
rect 2 21 5 41
rect 13 26 16 41
rect 24 33 26 41
rect 25 29 26 33
rect 13 22 14 26
rect 13 21 16 22
rect 24 21 26 29
rect 30 21 32 41
<< polycontact >>
rect 14 308 18 312
rect 21 301 25 305
rect 16 284 20 288
rect 16 264 20 268
rect 13 244 17 248
rect 17 226 21 230
rect 17 216 21 220
rect 16 209 20 213
rect 14 198 18 202
rect 14 153 18 157
rect 17 142 21 146
rect 17 135 21 139
rect 13 117 17 121
rect 13 99 17 103
rect 18 78 22 82
rect 16 66 20 70
rect 16 46 20 50
rect 21 29 25 33
rect 14 22 18 26
<< metal1 >>
rect 2 323 5 327
rect 30 323 32 327
rect 2 314 5 318
rect 30 314 32 318
rect 18 308 32 311
rect 2 302 21 305
rect 13 278 25 281
rect 9 271 16 274
rect 20 271 25 274
rect 2 262 5 266
rect 30 262 32 266
rect -3 251 -2 254
rect 2 250 5 254
rect 9 251 36 254
rect 9 237 23 240
rect -3 230 17 233
rect 21 230 36 233
rect -3 216 5 219
rect 9 216 17 219
rect 21 216 36 219
rect 2 197 5 201
rect 14 178 18 198
rect 30 197 32 201
rect -3 175 25 178
rect 29 175 36 178
rect -3 168 32 172
rect -3 161 25 164
rect 29 161 36 164
rect 2 154 5 158
rect 14 157 18 161
rect 30 154 32 158
rect 21 142 25 146
rect -3 136 5 139
rect 9 136 17 139
rect 21 136 36 139
rect -3 114 13 117
rect 17 114 36 117
rect 9 107 23 110
rect -3 92 -2 96
rect 2 93 5 96
rect 9 93 36 96
rect 2 92 36 93
rect 5 86 17 89
rect 21 86 29 89
rect -3 78 18 79
rect 22 78 36 79
rect -3 76 36 78
rect 2 68 5 72
rect 30 68 32 72
rect 9 60 16 63
rect 20 60 25 63
rect 13 53 25 56
rect 2 29 21 32
rect 18 23 32 26
rect 2 16 5 20
rect 30 16 32 20
rect -2 4 5 8
rect 30 4 32 8
<< m2contact >>
rect 5 334 9 338
rect -2 323 2 327
rect 32 323 36 327
rect -2 314 2 318
rect 32 314 36 318
rect 32 307 36 311
rect -2 301 2 305
rect 16 288 20 292
rect 9 278 13 282
rect 16 271 20 275
rect -2 262 2 266
rect 12 264 16 268
rect 32 262 36 266
rect -2 250 2 254
rect 17 244 21 248
rect 5 236 9 240
rect 17 230 21 234
rect 9 223 13 227
rect 5 215 9 219
rect 12 209 16 213
rect -2 197 2 201
rect 32 197 36 201
rect 25 175 29 179
rect 32 168 36 172
rect 25 161 29 165
rect -2 154 2 158
rect 32 154 36 158
rect 25 142 29 146
rect 5 136 9 140
rect 5 124 9 128
rect 13 113 17 117
rect 5 107 9 111
rect 17 99 21 103
rect -2 92 2 96
rect 17 85 21 89
rect -2 68 2 72
rect 12 66 16 70
rect 32 68 36 72
rect 16 59 20 63
rect 9 52 13 56
rect 16 42 20 46
rect -2 29 2 33
rect 32 23 36 27
rect -2 16 2 20
rect 32 16 36 20
rect -2 8 2 12
rect 32 4 36 8
<< metal2 >>
rect 5 338 8 344
rect 15 338 18 344
rect 9 334 10 338
rect -2 327 2 334
rect -2 318 2 323
rect 15 323 18 334
rect 32 327 36 344
rect 15 320 19 323
rect -2 305 2 314
rect -2 266 2 301
rect 16 296 19 320
rect 32 318 36 323
rect 32 311 36 314
rect 16 292 20 296
rect -2 254 2 262
rect -2 201 2 250
rect 9 227 12 278
rect 16 275 19 288
rect 32 266 36 307
rect 21 244 28 248
rect 21 230 22 234
rect -2 158 2 197
rect -2 96 2 154
rect 5 140 8 215
rect 19 197 22 230
rect 13 194 22 197
rect 5 111 9 124
rect 13 117 16 194
rect 25 185 28 244
rect 19 182 28 185
rect 32 201 36 262
rect 19 139 22 182
rect 25 165 29 175
rect 32 172 36 197
rect 32 158 36 168
rect 19 136 23 139
rect -2 72 2 92
rect -2 33 2 68
rect 9 56 12 110
rect 20 103 23 136
rect 21 99 23 103
rect 17 89 21 99
rect 26 86 29 142
rect 24 82 29 86
rect 16 46 19 59
rect 9 42 16 46
rect -2 20 2 29
rect -2 12 2 16
rect 24 15 28 82
rect 5 0 8 12
rect 13 11 28 15
rect 32 72 36 154
rect 32 27 36 68
rect 32 20 36 23
rect 13 7 17 11
rect 13 0 17 3
rect 32 8 36 16
rect 32 0 36 4
<< m3contact >>
rect 15 334 19 338
rect 5 330 9 334
rect 12 205 16 209
rect 5 42 9 46
rect 5 12 9 16
rect 13 3 17 7
<< metal3 >>
rect 4 334 10 344
rect 4 330 5 334
rect 9 330 10 334
rect 4 327 10 330
rect 14 338 20 344
rect 14 334 15 338
rect 19 334 20 338
rect 14 327 20 334
rect 3 322 10 327
rect 3 48 8 322
rect 11 209 17 210
rect 11 205 12 209
rect 16 205 17 209
rect 11 204 17 205
rect 11 56 16 204
rect 11 51 18 56
rect 3 46 10 48
rect 3 42 5 46
rect 9 42 10 46
rect 3 41 10 42
rect 13 21 18 51
rect 3 16 18 21
rect 3 12 5 16
rect 9 12 10 16
rect 3 11 10 12
rect 3 0 8 11
rect 12 7 18 8
rect 12 3 13 7
rect 17 3 18 7
rect 12 2 18 3
rect 12 0 17 2
<< m3p >>
rect 0 0 34 344
<< labels >>
rlabel metal1 -3 76 -3 76 1 reset
rlabel metal1 -3 168 -3 168 3 gnd
rlabel metal1 -3 175 -3 175 5 en2_S
rlabel metal1 -3 92 -3 92 1 vdd
rlabel metal1 -3 114 -3 114 5 S
rlabel metal1 -3 216 -3 216 1 en1_S
rlabel metal3 14 344 14 344 5 Q
rlabel metal3 5 1 5 1 1 bm_in
rlabel metal3 12 0 12 0 1 D
rlabel metal3 4 344 4 344 5 bm_out
<< end >>
