
.SUBCKT power_gate_cell sleep vvdd vdd
M0 vvdd sleep vdd vdd p l=0.6u w=7.5u m=3
.ENDS power_gate_cell
