magic
tech scmos
timestamp 1614203569
<< nwell >>
rect -2 89 17 173
rect -2 0 19 89
<< pwell >>
rect 17 89 36 173
rect 19 0 36 89
<< ntransistor >>
rect 23 140 30 142
rect 23 131 30 133
rect 23 122 30 124
rect 23 114 30 116
rect 26 76 30 78
rect 26 62 30 64
rect 26 44 30 48
rect 26 18 30 38
<< ptransistor >>
rect 5 140 11 142
rect 5 122 11 124
rect 5 97 11 99
rect 5 76 13 78
rect 5 62 13 64
rect 5 44 13 48
rect 5 18 13 38
<< ndiffusion >>
rect 23 143 26 147
rect 23 142 30 143
rect 23 133 30 140
rect 23 124 30 131
rect 23 116 30 122
rect 23 107 30 114
rect 27 104 30 107
rect 29 79 30 83
rect 26 78 30 79
rect 26 69 30 76
rect 26 64 30 65
rect 26 61 30 62
rect 29 57 30 61
rect 29 49 30 53
rect 26 48 30 49
rect 26 43 30 44
rect 29 39 30 43
rect 26 38 30 39
rect 26 17 30 18
<< pdiffusion >>
rect 9 143 11 147
rect 5 142 11 143
rect 5 124 11 140
rect 5 121 11 122
rect 9 117 11 121
rect 9 100 11 104
rect 5 99 11 100
rect 5 94 11 97
rect 9 90 11 94
rect 9 79 13 83
rect 5 78 13 79
rect 5 69 13 76
rect 9 65 13 69
rect 5 64 13 65
rect 5 61 13 62
rect 9 57 13 61
rect 9 49 13 53
rect 5 48 13 49
rect 5 43 13 44
rect 9 39 13 43
rect 5 38 13 39
rect 5 17 13 18
rect 9 13 13 17
<< ndcontact >>
rect 26 143 30 147
rect 23 103 27 107
rect 25 79 29 83
rect 26 65 30 69
rect 25 57 29 61
rect 25 49 29 53
rect 25 39 29 43
rect 26 13 30 17
<< pdcontact >>
rect 5 143 9 147
rect 5 117 9 121
rect 5 100 9 104
rect 5 90 9 94
rect 5 79 9 83
rect 5 65 9 69
rect 5 57 9 61
rect 5 49 9 53
rect 5 39 9 43
rect 5 13 9 17
<< psubstratepcontact >>
rect 26 4 30 8
<< nsubstratencontact >>
rect 5 4 9 8
<< polysilicon >>
rect 3 140 5 142
rect 11 140 23 142
rect 30 140 32 142
rect 21 131 23 133
rect 30 131 32 133
rect 3 122 5 124
rect 11 122 23 124
rect 30 122 32 124
rect 21 114 23 116
rect 30 114 32 116
rect 3 97 5 99
rect 11 97 13 99
rect 3 76 5 78
rect 13 76 18 78
rect 22 76 26 78
rect 30 76 32 78
rect 3 62 5 64
rect 13 63 16 64
rect 20 63 26 64
rect 13 62 26 63
rect 30 62 32 64
rect 3 44 5 48
rect 13 47 26 48
rect 13 44 16 47
rect 20 44 26 47
rect 30 44 32 48
rect 2 18 5 38
rect 13 23 16 38
rect 24 30 26 38
rect 25 26 26 30
rect 13 19 14 23
rect 13 18 16 19
rect 24 18 26 26
rect 30 18 32 38
<< polycontact >>
rect 14 142 18 146
rect 17 131 21 135
rect 17 124 21 128
rect 17 114 21 118
rect 13 96 17 100
rect 18 75 22 79
rect 16 63 20 67
rect 16 43 20 47
rect 21 26 25 30
rect 14 19 18 23
<< metal1 >>
rect -3 156 32 160
rect -3 150 36 153
rect 2 143 5 147
rect 14 146 18 150
rect 30 143 32 147
rect -3 125 17 128
rect 21 125 36 128
rect -3 111 36 114
rect 9 104 23 107
rect -3 89 -2 93
rect 2 90 5 93
rect 9 90 36 93
rect 2 89 36 90
rect 5 83 17 86
rect 21 83 29 86
rect -3 75 18 76
rect 22 75 36 76
rect -3 73 36 75
rect 2 65 5 69
rect 30 65 32 69
rect 9 57 16 60
rect 20 57 25 60
rect 13 50 25 53
rect 2 26 21 29
rect 18 20 32 23
rect 2 13 5 17
rect 30 13 32 17
rect 2 4 5 8
rect 30 4 32 8
<< m2contact >>
rect 32 156 36 160
rect -2 143 2 147
rect 32 143 36 147
rect 21 131 25 135
rect 9 117 13 121
rect 5 104 9 108
rect 17 96 21 100
rect -2 89 2 93
rect 17 82 21 86
rect -2 65 2 69
rect 12 63 16 67
rect 32 65 36 69
rect 16 56 20 60
rect 9 49 13 53
rect 16 39 20 43
rect -2 26 2 30
rect 32 20 36 24
rect -2 13 2 17
rect 32 13 36 17
rect -2 4 2 8
rect 32 4 36 8
<< metal2 >>
rect 15 164 19 173
rect -2 147 2 163
rect 32 160 36 173
rect -2 93 2 143
rect 32 147 36 156
rect 25 131 28 135
rect -2 69 2 89
rect -2 30 2 65
rect 9 53 12 117
rect 17 86 21 96
rect 16 43 19 56
rect 10 39 16 43
rect 16 35 20 39
rect -2 17 2 26
rect -2 8 2 13
rect 24 9 28 131
rect -2 0 2 4
rect 13 6 28 9
rect 32 69 36 143
rect 32 24 36 65
rect 32 17 36 20
rect 32 8 36 13
rect 13 0 17 2
rect 32 0 36 4
<< m3contact >>
rect 15 160 19 164
rect 6 39 10 43
rect 13 2 17 6
<< metal3 >>
rect 14 164 20 173
rect 14 160 15 164
rect 19 160 20 164
rect 6 155 20 160
rect 6 49 11 155
rect 5 43 11 49
rect 5 39 6 43
rect 10 39 11 43
rect 5 38 11 39
rect 12 6 19 7
rect 12 2 13 6
rect 17 2 19 6
rect 12 0 19 2
<< m3p >>
rect 0 0 34 173
<< labels >>
rlabel metal1 -3 73 -3 73 1 reset
rlabel metal1 -3 150 -3 150 1 en2_S
rlabel metal1 -3 111 -3 111 1 S
rlabel metal1 -3 125 -3 125 1 en1_S
rlabel metal1 -3 89 -3 89 1 vdd
rlabel metal1 -3 156 -3 156 3 gnd
rlabel metal3 13 0 13 0 1 D
rlabel metal3 15 173 15 173 5 Q
<< end >>
