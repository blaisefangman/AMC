magic
tech scmos
timestamp 1615817584
<< nwell >>
rect 0 -2 44 40
<< ptransistor >>
rect 11 26 36 28
rect 11 18 36 20
rect 11 10 36 12
<< pdiffusion >>
rect 11 29 13 33
rect 19 29 23 33
rect 32 29 36 33
rect 11 28 36 29
rect 11 25 36 26
rect 11 21 17 25
rect 26 21 30 25
rect 11 20 36 21
rect 11 17 36 18
rect 11 13 13 17
rect 19 13 23 17
rect 32 13 36 17
rect 11 12 36 13
rect 11 9 36 10
rect 11 5 17 9
rect 26 5 30 9
<< pdcontact >>
rect 13 29 19 33
rect 23 29 32 33
rect 17 21 26 25
rect 30 21 36 25
rect 13 13 19 17
rect 23 13 32 17
rect 17 5 26 9
rect 30 5 36 9
<< nsubstratencontact >>
rect 3 31 7 35
<< polysilicon >>
rect 10 26 11 28
rect 36 26 38 28
rect 10 18 11 20
rect 36 18 38 20
rect 10 10 11 12
rect 36 10 38 12
<< polycontact >>
rect 6 24 10 28
rect 6 16 10 20
rect 6 8 10 12
<< metal1 >>
rect 0 36 19 40
rect 23 36 32 40
rect 36 36 44 40
rect 3 35 7 36
rect 6 20 10 24
rect 2 19 6 20
rect 0 16 6 19
rect 39 19 43 20
rect 6 12 10 16
rect 39 16 44 19
rect 0 -2 44 2
<< m2contact >>
rect 19 36 23 40
rect 32 36 36 40
rect 19 29 23 33
rect 32 29 36 33
rect 2 20 6 24
rect 13 21 17 25
rect 26 21 30 25
rect 39 20 43 24
rect 19 13 23 17
rect 32 13 36 17
rect 13 5 17 9
rect 26 5 30 9
<< metal2 >>
rect 13 25 16 40
rect 20 33 23 36
rect 13 9 16 21
rect 20 17 23 29
rect 13 -2 16 5
rect 20 -2 23 13
rect 26 25 29 40
rect 33 33 36 36
rect 26 9 29 21
rect 33 17 36 29
rect 26 -2 29 5
rect 33 -2 36 13
<< m3contact >>
rect 2 16 6 20
rect 39 16 43 20
<< metal3 >>
rect 0 20 44 21
rect 0 16 2 20
rect 6 16 39 20
rect 43 16 44 20
rect 0 15 44 16
<< m3p >>
rect 0 0 44 38
<< labels >>
rlabel metal1 0 16 0 16 3 sleep
rlabel metal2 13 -2 13 -2 1 vvdd
rlabel metal2 20 -2 20 -2 1 vdd
rlabel metal2 26 -2 26 -2 1 vvdd
rlabel metal2 33 -2 33 -2 1 vdd
<< end >>
