magic
tech scmos
timestamp 1615755140
<< nwell >>
rect 37 -2 79 68
rect 137 -2 166 68
<< pwell >>
rect 0 -2 37 68
rect 79 -2 137 68
<< ntransistor >>
rect 91 48 95 50
rect 121 48 125 50
rect 27 39 31 41
rect 121 40 125 42
rect 27 31 31 33
rect 91 32 95 34
rect 121 32 125 34
rect 91 24 95 26
rect 91 16 95 18
rect 121 16 125 18
<< ptransistor >>
rect 69 48 73 50
rect 143 48 147 50
rect 44 39 52 41
rect 143 40 147 42
rect 44 31 52 33
rect 69 32 73 34
rect 143 32 147 34
rect 69 24 73 26
rect 69 16 73 18
rect 143 16 147 18
<< ndiffusion >>
rect 91 50 95 51
rect 121 50 125 51
rect 27 41 31 42
rect 91 47 95 48
rect 121 47 125 48
rect 121 42 125 43
rect 27 38 31 39
rect 27 33 31 34
rect 121 39 125 40
rect 91 34 95 35
rect 121 34 125 35
rect 27 30 31 31
rect 91 31 95 32
rect 121 31 125 32
rect 91 26 95 27
rect 91 23 95 24
rect 91 18 95 19
rect 121 18 125 19
rect 91 15 95 16
rect 121 15 125 16
<< pdiffusion >>
rect 69 50 73 51
rect 143 50 147 51
rect 44 42 48 46
rect 44 41 52 42
rect 69 47 73 48
rect 143 47 147 48
rect 143 42 147 43
rect 44 38 52 39
rect 44 34 48 38
rect 69 34 73 35
rect 44 33 52 34
rect 143 39 147 40
rect 143 34 147 35
rect 69 31 73 32
rect 44 30 52 31
rect 44 26 48 30
rect 69 26 73 27
rect 143 31 147 32
rect 69 23 73 24
rect 69 18 73 19
rect 143 18 147 19
rect 69 15 73 16
rect 143 15 147 16
<< ndcontact >>
rect 91 51 95 55
rect 121 51 125 55
rect 27 42 31 46
rect 91 43 95 47
rect 121 43 125 47
rect 27 34 31 38
rect 91 35 95 39
rect 121 35 125 39
rect 27 26 31 30
rect 91 27 95 31
rect 121 27 125 31
rect 91 19 95 23
rect 121 19 125 23
rect 91 11 95 15
rect 121 11 125 15
<< pdcontact >>
rect 69 51 73 55
rect 143 51 147 55
rect 48 42 52 46
rect 69 43 73 47
rect 143 43 147 47
rect 48 34 52 38
rect 69 35 73 39
rect 143 35 147 39
rect 48 26 52 30
rect 69 27 73 31
rect 143 27 147 31
rect 69 19 73 23
rect 143 19 147 23
rect 69 11 73 15
rect 143 11 147 15
<< psubstratepcontact >>
rect 105 32 109 36
rect 22 5 26 9
<< nsubstratencontact >>
rect 52 6 56 10
rect 157 8 161 12
<< polysilicon >>
rect 63 48 69 50
rect 73 48 75 50
rect 89 48 91 50
rect 95 48 98 50
rect 102 48 121 50
rect 125 48 127 50
rect 141 48 143 50
rect 147 48 154 50
rect 63 44 65 48
rect 24 39 27 41
rect 31 39 44 41
rect 52 40 61 41
rect 52 39 65 40
rect 118 40 121 42
rect 125 40 143 42
rect 147 41 154 42
rect 147 40 150 41
rect 20 31 27 33
rect 31 31 33 33
rect 38 31 44 33
rect 52 31 54 33
rect 67 32 69 34
rect 73 32 91 34
rect 95 32 97 34
rect 119 32 121 34
rect 125 32 143 34
rect 147 32 149 34
rect 66 24 69 26
rect 73 24 91 26
rect 95 24 98 26
rect 66 16 69 18
rect 73 16 75 18
rect 89 16 91 18
rect 95 16 121 18
rect 125 16 127 18
rect 141 16 143 18
rect 147 16 150 18
<< polycontact >>
rect 98 48 102 52
rect 150 50 154 54
rect 61 40 65 44
rect 80 34 84 38
rect 114 38 118 42
rect 150 37 154 41
rect 20 27 24 31
rect 38 27 42 31
rect 62 24 66 28
rect 98 24 102 28
rect 132 28 136 32
rect 112 18 116 22
rect 62 14 66 18
rect 150 16 154 20
<< metal1 >>
rect 0 64 42 68
rect 46 64 69 68
rect 73 64 143 68
rect 147 64 166 68
rect 0 58 61 61
rect 65 58 112 61
rect 116 58 166 61
rect 0 51 69 54
rect 73 51 91 55
rect 125 51 132 55
rect 136 51 143 55
rect 150 54 154 58
rect 161 51 166 54
rect 31 42 48 45
rect 52 42 58 45
rect 0 27 20 31
rect 27 23 31 26
rect 48 23 52 26
rect 27 20 52 23
rect 0 13 34 17
rect 55 18 58 42
rect 73 43 91 47
rect 125 43 143 47
rect 147 44 166 47
rect 80 42 84 43
rect 62 35 69 37
rect 62 34 73 35
rect 95 35 102 39
rect 62 28 66 34
rect 98 28 102 35
rect 114 32 118 38
rect 114 31 125 32
rect 114 29 121 31
rect 150 31 154 37
rect 73 19 91 23
rect 55 14 62 18
rect 98 15 102 24
rect 147 27 154 31
rect 132 23 136 24
rect 125 19 143 23
rect 62 8 66 14
rect 73 11 80 15
rect 84 11 91 15
rect 98 12 121 15
rect 125 11 143 15
rect 62 5 98 8
rect 150 8 153 16
rect 102 5 153 8
rect 22 2 26 5
rect 0 -2 27 2
rect 31 -2 91 2
rect 95 -2 105 2
rect 109 -2 121 2
rect 125 -2 166 2
<< m2contact >>
rect 42 64 46 68
rect 69 64 73 68
rect 143 64 147 68
rect 61 57 65 61
rect 112 57 116 61
rect 132 51 136 55
rect 157 50 161 54
rect 23 35 27 39
rect 44 34 48 38
rect 34 27 38 31
rect 34 13 38 17
rect 48 16 52 20
rect 61 44 65 48
rect 98 44 102 48
rect 80 38 84 42
rect 73 27 77 31
rect 87 27 91 31
rect 105 28 109 32
rect 125 35 129 39
rect 139 35 143 39
rect 154 37 158 41
rect 112 22 116 26
rect 132 24 136 28
rect 48 6 52 10
rect 80 11 84 15
rect 98 5 102 9
rect 157 12 161 16
rect 27 -2 31 2
rect 91 -2 95 2
rect 105 -2 109 2
rect 121 -2 125 2
<< metal2 >>
rect 27 2 31 39
rect 42 38 46 64
rect 61 48 65 57
rect 42 34 44 38
rect 34 17 37 27
rect 42 10 45 34
rect 52 16 55 46
rect 69 27 73 64
rect 98 48 102 52
rect 80 15 84 38
rect 42 6 48 10
rect 91 2 95 31
rect 98 9 102 44
rect 105 2 109 28
rect 112 26 116 57
rect 121 2 125 39
rect 132 28 136 51
rect 143 16 147 64
rect 154 50 157 54
rect 161 51 166 54
rect 154 41 158 46
rect 143 12 157 16
<< m3contact >>
rect 52 46 56 50
rect 154 46 158 50
<< metal3 >>
rect 51 50 57 51
rect 153 50 161 51
rect 51 46 52 50
rect 56 46 154 50
rect 158 46 161 50
rect 51 45 161 46
<< m3p >>
rect 0 0 166 66
<< labels >>
rlabel metal1 166 51 166 51 7 out
rlabel metal1 166 44 166 44 7 out_bar
rlabel metal1 0 58 0 58 3 clk
rlabel metal1 0 66 0 66 4 vdd
rlabel metal1 0 51 0 51 3 in
rlabel metal1 0 27 0 27 3 rst0
rlabel metal1 0 13 0 13 3 rst1
rlabel metal1 0 0 0 0 2 gnd
<< end >>
