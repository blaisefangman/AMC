magic
tech scmos
timestamp 1614182919
<< nwell >>
rect -6 128 34 273
rect -6 51 34 83
<< pwell >>
rect -6 273 34 330
rect -6 83 34 128
rect -6 28 34 51
<< ntransistor >>
rect 12 301 14 319
rect 12 279 14 288
rect 20 279 22 288
rect 9 118 11 122
rect 17 118 19 122
rect 13 37 15 45
rect 21 37 23 45
<< ptransistor >>
rect 12 249 14 267
rect 20 249 22 267
rect 10 199 12 223
rect 21 168 23 192
rect 9 134 11 142
rect 17 134 19 142
rect 13 57 15 65
rect 21 57 23 65
<< ndiffusion >>
rect 11 301 12 319
rect 14 301 15 319
rect 11 279 12 288
rect 14 279 15 288
rect 19 279 20 288
rect 22 279 23 288
rect 8 118 9 122
rect 11 118 12 122
rect 16 118 17 122
rect 19 118 20 122
rect 12 37 13 45
rect 15 37 16 45
rect 20 37 21 45
rect 23 37 24 45
<< pdiffusion >>
rect 7 265 12 267
rect 11 251 12 265
rect 7 249 12 251
rect 14 265 20 267
rect 14 251 15 265
rect 19 251 20 265
rect 14 249 20 251
rect 22 265 27 267
rect 22 251 23 265
rect 22 249 27 251
rect 9 199 10 223
rect 12 199 13 223
rect 20 181 21 192
rect 16 168 21 181
rect 23 168 24 192
rect 8 134 9 142
rect 11 134 12 142
rect 16 134 17 142
rect 19 134 20 142
rect 8 63 13 65
rect 12 59 13 63
rect 8 57 13 59
rect 15 63 21 65
rect 15 59 16 63
rect 20 59 21 63
rect 15 57 21 59
rect 23 63 28 65
rect 23 59 24 63
rect 23 57 28 59
<< ndcontact >>
rect 7 301 11 319
rect 15 301 19 319
rect 7 279 11 288
rect 15 279 19 288
rect 23 279 27 288
rect 4 118 8 122
rect 12 118 16 122
rect 20 118 24 122
rect 8 37 12 45
rect 16 37 20 45
rect 24 37 28 45
<< pdcontact >>
rect 7 251 11 265
rect 15 251 19 265
rect 23 251 27 265
rect 5 199 9 223
rect 13 199 17 223
rect 16 181 20 192
rect 24 168 28 192
rect 4 134 8 142
rect 12 134 16 142
rect 20 134 24 142
rect 8 59 12 63
rect 16 59 20 63
rect 24 59 28 63
<< psubstratepcontact >>
rect -2 318 2 322
rect 16 104 20 108
rect -2 37 2 41
<< nsubstratencontact >>
rect 12 233 16 237
rect 12 156 16 160
rect 27 69 31 73
<< polysilicon >>
rect 12 319 14 321
rect 12 300 14 301
rect 12 298 31 300
rect 3 293 22 295
rect 3 276 5 293
rect 12 288 14 290
rect 20 288 22 293
rect 3 272 4 276
rect 3 230 5 272
rect 12 267 14 279
rect 20 267 22 279
rect 12 244 14 249
rect 20 247 22 249
rect 12 242 22 244
rect 23 226 25 240
rect 10 223 12 225
rect 10 167 12 199
rect 29 195 31 298
rect 21 193 31 195
rect 21 192 23 193
rect 21 167 23 168
rect 10 165 27 167
rect 5 149 7 160
rect 25 153 27 165
rect 5 147 31 149
rect 9 142 11 144
rect 17 142 19 144
rect 9 122 11 134
rect 17 131 19 134
rect 18 127 19 131
rect 17 122 19 127
rect 4 100 6 111
rect 4 85 6 96
rect 9 92 11 118
rect 17 116 19 118
rect 4 83 15 85
rect 29 83 31 147
rect 13 65 15 79
rect 21 79 27 81
rect 21 65 23 79
rect 13 55 15 57
rect 6 49 15 51
rect 13 45 15 49
rect 21 45 23 57
rect 13 35 15 37
rect 21 30 23 37
rect 6 28 23 30
<< polycontact >>
rect 4 272 8 276
rect 22 240 26 244
rect 3 226 7 230
rect 21 222 25 226
rect 3 160 7 164
rect 21 153 25 157
rect 14 127 18 131
rect 2 111 6 115
rect 2 96 6 100
rect 9 88 13 92
rect 11 79 15 83
rect 27 79 31 83
rect 2 49 6 53
rect 2 28 6 32
<< metal1 >>
rect 2 322 34 326
rect 7 319 11 322
rect 15 288 18 301
rect 7 276 11 279
rect 8 272 11 276
rect 7 265 11 272
rect 7 249 11 251
rect 15 265 19 267
rect 23 265 27 279
rect 15 246 18 251
rect 13 243 18 246
rect 23 244 27 251
rect 13 237 16 243
rect 26 240 27 244
rect 0 233 12 237
rect 16 233 27 237
rect 31 233 34 237
rect 3 223 7 226
rect 3 199 5 223
rect 3 164 6 199
rect 25 192 28 225
rect 18 169 24 173
rect 12 160 27 164
rect 12 142 16 156
rect 21 142 24 153
rect 4 131 8 134
rect 4 127 14 131
rect 4 122 8 127
rect 21 122 24 134
rect 4 115 8 118
rect 6 111 8 115
rect 12 108 16 118
rect 2 104 16 108
rect -2 88 9 91
rect 13 88 34 91
rect 2 53 5 88
rect 25 65 27 69
rect 25 63 28 65
rect 9 45 12 59
rect 16 45 20 59
rect 25 45 27 48
rect 12 37 13 45
rect 9 36 13 37
rect 10 32 13 36
rect 10 28 27 32
rect 2 25 6 28
<< m2contact >>
rect -2 322 2 326
rect 27 233 31 237
rect 13 223 17 227
rect 17 192 21 196
rect 14 169 18 173
rect 27 160 31 164
rect -2 104 2 108
rect 27 65 31 69
rect 27 45 31 49
rect -2 41 2 45
rect 27 28 31 32
rect 2 21 6 25
<< metal2 >>
rect -2 326 2 330
rect -2 108 2 322
rect 9 319 14 330
rect 10 227 14 319
rect 10 223 13 227
rect 10 202 14 223
rect 8 199 14 202
rect 8 149 11 199
rect 20 196 24 330
rect 8 146 12 149
rect -2 45 2 104
rect -2 37 2 41
rect -2 33 -1 37
rect 2 0 5 21
rect 9 0 12 146
rect 15 0 18 169
rect 21 21 24 196
rect 27 237 31 330
rect 27 164 31 233
rect 27 69 31 160
rect 21 18 25 21
rect 22 0 25 18
rect 28 0 31 24
<< m3contact >>
rect -1 33 3 37
rect 27 49 31 53
rect 27 24 31 28
<< metal3 >>
rect 26 53 32 54
rect 26 49 27 53
rect 31 49 32 53
rect 26 38 32 49
rect -2 37 32 38
rect -2 33 -1 37
rect 3 33 32 37
rect -2 32 4 33
rect 24 28 32 29
rect 24 24 27 28
rect 31 24 32 28
rect 24 23 32 24
rect 24 0 29 23
<< m3p >>
rect 0 0 34 330
<< labels >>
flabel metal1 34 233 34 233 6 FreeSans 26 180 0 0 vdd
flabel metal1 34 322 34 322 6 FreeSans 26 180 0 0 gnd
flabel metal1 34 88 34 88 6 FreeSans 26 180 0 0 en
rlabel metal2 20 330 20 330 5 bl
rlabel metal2 9 330 9 330 5 br
rlabel metal2 15 1 15 1 1 dout1
rlabel metal2 2 1 2 1 1 dout_bar
rlabel metal3 24 0 24 0 1 dout
<< properties >>
string path 270.000 468.000 270.000 486.000 288.000 486.000 288.000 468.000 270.000 468.000 
<< end >>
